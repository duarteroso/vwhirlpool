module vwhirlpool
